Library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

entity FREQ_DEVIDER is
	port(CLK:in STD_LOGIC;
		  CLK1HZ,CLK2HZ,CLK390KHZ:out STD_LOGIC);
end FREQ_DEVIDER;

architecture Behaviorual of FREQ_DEVIDER is
	COMPONENT DIVCLKTO1HZ
	port(MCLK:in STD_LOGIC;
	     CLK1HZ:out STD_LOGIC);
	end COMPONENT;
	
	COMPONENT DIVCLKTO2HZ
	port(MCLK:in STD_LOGIC;
	     CLK2HZ:out STD_LOGIC);
	end COMPONENT;
	
	COMPONENT DIVCLKTO390KHZ
	port(MCLK:in STD_LOGIC;
	     CLK390KHZ:out STD_LOGIC);
	end COMPONENT;
	begin
	GENCLK1HZ:DIVCLKTO1HZ port map(CLK,CLK1HZ);
	GENCLK2HZ:DIVCLKTO2HZ port map(CLK,CLK2HZ);
	GENCLK390KHZ:DIVCLKTO390KHZ port map(CLK,CLK390KHZ);
end Behaviorual;